`define N 5'b10011